* 3x3 Resistor Grid Netlist
* simple test for Cholesky factorization

*.options METHOD=tr
*.tran 0.5 2.6

*.options iter spd
* passive elementsns
*.options sparse
*.options


R00 _n_00_00_  _n_25_00_  4
R01 _n_25_00_  _n_50_00_  32

R02 _n_00_00_  _n_00_25_  18
R03 _n_25_00_  _n_25_25_  15
R04 _n_50_00_  _n_50_25_  92

R05 _n_00_25_  _n_25_25_  15
R06 _n_25_25_  _n_50_25_  28

R07 _n_00_25_  _n_00_50_  33
R08 _n_25_25_  _n_25_50_  29
R09 _n_50_25_  _n_50_50_  12

R10 _n_00_50_  _n_25_50_  48
R11 _n_25_50_  _n_50_50_  90

C12 _n_25_50_ _n_00_50_ 10 

Rg1  _n_25_00_ 0 100
Rg2  _n_50_00_ 0 100

* current source
Isrc _n_00_00_  0 10 exp (10 5 1 0.2 2 0.5)


* options setup
.options spd iter


* required simulation
 .dc Isrc 0 10 0.1 
 *.dc Ia 0 10 0.1

* required output
.plot V(_n_00_00_) V(_n_00_50_)

.end
